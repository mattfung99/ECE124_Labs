    Mac OS X            	   2         �                                      ATTR       �   �                     �     com.apple.quarantine q/0082;5a6627a5;Outlook; 