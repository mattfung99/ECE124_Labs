    Mac OS X            	   2       C                                      ATTR      C   �   S                  �     com.apple.lastuseddate#PS          *  $com.apple.metadata:_kMDItemUserTags    *     com.apple.quarantine H�Z    Q2    bplist00�                            	q/0082;5aa005e5;Outlook; 